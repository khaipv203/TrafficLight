module display(
   input [5:0] bin,
   output [13:0] display
   );
   
    assign display = (bin == 6'b000000) ? 14'b00000010000001: //0
                (bin == 6'b000001) ? 14'b00000011001111: //1
                (bin == 6'b000010) ? 14'b00000010010010: //2
                (bin == 6'b000011) ? 14'b00000010000110: //3
                (bin == 6'b000100) ? 14'b00000011001100: //4
                (bin == 6'b000101) ? 14'b00000010100100: //5
                (bin == 6'b000110) ? 14'b00000010100000: //6
                (bin == 6'b000111) ? 14'b00000010001111: //7
                (bin == 6'b001000) ? 14'b00000010000000: //8
                (bin == 6'b001001) ? 14'b00000010000100: //9
                (bin == 6'b001010) ? 14'b00000010000001: //10
                (bin == 6'b001011) ? 14'b00000011001111: //11
                (bin == 6'b001100) ? 14'b00000010010010: //12
                (bin == 6'b001101) ? 14'b00000010000110: //13
                (bin == 6'b001110) ? 14'b00000011001100: //14
                (bin == 6'b001110) ? 14'b00000010100100: //15
                (bin == 6'b001111) ? 14'b00000010100000: //16
                (bin == 6'b010000) ? 14'b00000010001111: //17
                (bin == 6'b010001) ? 14'b00000010000000: //18
                (bin == 6'b010010) ? 14'b00000010000100: //19
                (bin == 6'b010011) ? 14'b00100100000001: //20
                (bin == 6'b010100) ? 14'b00100101001111: //21
                (bin == 6'b010101) ? 14'b00100100010010: //22
                (bin == 6'b010110) ? 14'b00100100000110: //23
                (bin == 6'b010111) ? 14'b00100101001100: //24
                (bin == 6'b011000) ? 14'b00100100100100: //25
                (bin == 6'b011001) ? 14'b00100100100000: //26
                (bin == 6'b011010) ? 14'b00100100001111: //27
                (bin == 6'b011011) ? 14'b00100100000000: //28
                (bin == 6'b011100) ? 14'b00100100000100: //29
                (bin == 6'b011101) ? 14'b00001100000001: //30
                (bin == 6'b011110) ? 14'b00001101001111: //31
                (bin == 6'b011111) ? 14'b00001100010010: //32
                (bin == 6'b100000) ? 14'b00001100000110: //33
                (bin == 6'b100001) ? 14'b00001101001100: //34
                (bin == 6'b100010) ? 14'b00001100100100: //35
                (bin == 6'b100011) ? 14'b00001100100000: //36
                (bin == 6'b100100) ? 14'b00001100001111: //37
                (bin == 6'b100101) ? 14'b00001100000000: //38
                (bin == 6'b100110) ? 14'b00001100000100: //39
                (bin == 6'b100111) ? 14'b10011000000001: //40
                (bin == 6'b101000) ? 14'b10011001001111: //41
                (bin == 6'b101001) ? 14'b10011000010010: //42
                (bin == 6'b101010) ? 14'b10011000000110: //43
                (bin == 6'b101011) ? 14'b10011001001100: //44
                (bin == 6'b101100) ? 14'b10011000100100: //45
                (bin == 6'b101101) ? 14'b10011000100000: //46
                (bin == 6'b101110) ? 14'b10011000001111: //47
                (bin == 6'b101111) ? 14'b10011000000000: //48
                (bin == 6'b110000) ? 14'b10011000000100: //49
                (bin == 6'b110001) ? 14'b01001000000001: //50
                (bin == 6'b110010) ? 14'b01001001001111: //51
                (bin == 6'b110011) ? 14'b01001000010010: //52
                (bin == 6'b110100) ? 14'b01001000000110: //53
                (bin == 6'b110101) ? 14'b01001001001100: //54
                (bin == 6'b110110) ? 14'b01001000100100: //55
                (bin == 6'b110111) ? 14'b01001000100000: //56
                (bin == 6'b111000) ? 14'b01001000001111: //57
                (bin == 6'b111001) ? 14'b01001000000000: //58
                (bin == 6'b111010) ? 14'b01001000000100: 14'b11111111111111; //59

endmodule